module LAB2_MUX(SW,KEY,LEDR);
	input [9:0] SW;
	input [3:0] KEY;
	output [9:0] LEDR;
	
	//lab2_1 zad1(SW, LEDR);
	//lab2_2 zad2({KEY[0], KEY[1], KEY[2], KEY[3]}, {LEDR[0], LEDR[1], LEDR[2], LEDR[3]});
	lab2_3 zad3(SW, KEY, LEDR);
	
	// lab2_4 zad4(SW,LEDR,KEY); 
 	
	
	
	//lab2_5 zad5(SW,KEY,LEDR);
	//lab2_6 zad6();
	//lab2_7 zad7();
	//lab2_8 zad8();
	//lab2_9 zad9();
	//lab2_10 zad10();
	//lab2_11 zad11();
	//lab2_12 zad12();
endmodule